Vin 0 1 5
X 1 2 SK1
X 2 3 NIA
Vout 3
.end