R1 1 2 1k
R2 2 0 1k
.declare_subckt 1 2
.end
