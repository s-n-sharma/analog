R1 1 2 1k
X 2 3 RC
.declare_subckt 1 3
.end 