Vin 0 1 5
X 1 2 RC
IOP 2 3 3
.end 
