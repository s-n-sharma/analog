R1 1 2 1k
R2 2 3 1k 
IOP 3 4 4 
C1 2 4 1u
C2 3 0 1u
.declare_subckt 1 4 
.end
