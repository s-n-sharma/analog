R1 1 2 1k
C1 2 0 1u
.declare_subckt 1 2
.ends