IOP 2 1 2
R1 2 3 1k
R2 3 0 1k
.declare_subckt 1 3
.end