Vin 0 1 5
X 1 2 RC
X 2 3 RC2
VOUT 3
.end
