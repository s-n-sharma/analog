IOP 1 2 3 
R2 2 0 1k 
R1 2 3 5k 
.declare_subckt 1 3 
.end